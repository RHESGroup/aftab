LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;


entity aftab_mem_controller is 
	
	PORT (

	);
end aftab_mem_controller;



architecture behv of aftab_mem_controller is

begin
-- memory controller implementation 
    

end architecture;