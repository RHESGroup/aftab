LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;


entity aftab_mem_datapath is 
	
	PORT (

	);
end aftab_mem_datapath;



architecture behv of aftab_mem_datapath is

begin
-- memory datapath implementation 
    

end architecture;